package pa_Package;

  parameter PARAMETER   = 1;
  localparam PARAMETER2 = 2;


endpackage
module mymodule();
    reg a = 0;
    reg b = 0;
endmodule;

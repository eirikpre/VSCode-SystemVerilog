

module excluded #(
  parameter A
)(
  input a
);

endmodule
module mymodule();
    reg a = 0;
endmodule;

/*
module abc
*/

 /*
               module 123
 */

/* dog

      module
cat */

module cat #(
)(
      logic ck
);
      // Module body
endmodule

module abc #(
)(
      logic ck
);
      // Module body
endmodule


module 123 #(
)(
      logic ck
);
      // Module body
endmodule



// No error

/*module abc
*/

/*
moduleabc
*/

/*

            text module 123
*/

/*
module (  123
*/

/*
Module www
*/

/* dog
     module
*/
module mymodule();
    reg a = 0;
        reg b = 1;
endmodule;

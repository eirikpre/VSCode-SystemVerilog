module mymodule();
    reg a = 0;
    reg b = 0;
    reg c = 1;
    reg d = 1;
endmodule;

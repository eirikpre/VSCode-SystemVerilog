`define MYMACRO 0
module mymodule();
    reg a = `MYMACRO;
    reg b = `MYMACRO;
endmodule;

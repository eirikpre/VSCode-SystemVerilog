`define MYMACRO 0
module mymodule();
    reg a = 0;
endmodule;
